module renderengine

import mathengine {Vertex}
pub struct Box {
	
}