module audioengine
/*
import os

pub fn play_sound(file str){
	if os.name == "nt"{
		os.system("start " + file)
	}else{
		os.system("afplay " + file)
	}
}
*/

pub fn play_sound(file string) {
	//os.system("afplay " + file)
}